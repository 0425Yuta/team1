module ALU(
	input wire clock,
	input wire[15:0] address_ram,
	input wire[15:0] q_ram,
	input wire[15:0] data_ram,
	input wire[15:0] address_rom,
	input wire[15:0] q_rom
);
endmodule
